library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity datapath_testbench is
--  Port ( );
end datapath_testbench;

architecture Behavioral of datapath_testbench is

begin


end Behavioral;
